--Copyright (C)2014-2025 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.11.03 (64-bit)
--Part Number: GW2A-LV18PG256C8/I7
--Device: GW2A-18
--Device Version: C
--Created Time: Sat Aug 30 21:22:18 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(0 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(12 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= gw_gnd & ad(12 downto 0);
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_08 => X"006C6CFE6CFE6C6C0000000000006C6C00300030307878300000000000000000",
            INIT_RAM_09 => X"0000000000060C0C00DC6676DC386C3800C6CC183066C60000183E603C067C18",
            INIT_RAM_0A => X"000018187E1818000000CC79FE78CC00000C18303030180C0030180C0C0C1830",
            INIT_RAM_0B => X"0002060C183060C00018180000000000000000007E0000000C18180000000000",
            INIT_RAM_0C => X"003C66603860663C007E660C3860663C007E181818181C18007CCEDEF6E6C67C",
            INIT_RAM_0D => X"001818183060667E003C66663E060C38003C6660603E067E00F060FE666C7870",
            INIT_RAM_0E => X"0C181800001818000018180000181800001C30607C66663C003C66663C66663C",
            INIT_RAM_0F => X"001800183060663C000C18306030180C00007E00007E00000030180C060C1830",
            INIT_RAM_10 => X"0078CC060606CC78007ECCCC7CCCCC7E0066667E66663C18003C06F6F6F6C67C",
            INIT_RAM_11 => X"00F8CCE60606CC78001E0C2C3C2C8CFE00FE8C2C3C2C8CFE003E6CCCCCCC6C3E",
            INIT_RAM_12 => X"00CECC6C3C6CCCCE003C6666606060F0003C18181818183C006666667E666666",
            INIT_RAM_13 => X"00386CC6C6C66C3800C6C6E6F6DECEC600C6C6D6FEFEEEC600FECC8C0C0C0C1E",
            INIT_RAM_14 => X"003C66701C0E663C00CECC6C7CCCCC7E00703C766666663C001E0C0C7CCCCC7E",
            INIT_RAM_15 => X"00C6EEFED6C6C6C600183C6666666666007E666666666666003C181818185A7E",
            INIT_RAM_16 => X"003C0C0C0C0C0C3C00FECC983062C6FE003C18183C66666600C66C38386CC6C6",
            INIT_RAM_17 => X"FE0000000000000000000000C66C3810003C30303030303C0080C06030180C06",
            INIT_RAM_18 => X"003C6606663C00000076CCCC7C0C0C0E00DC667C603C00000000000000301819",
            INIT_RAM_19 => X"3E607C6666DC0000001E0C0C1E0C6C38003C067E663C000000DC66667C606070",
            INIT_RAM_1A => X"00CE6C3C6CCC0C0E3C66666060600060003C1818181C001800CECCCCDC6C0C0E",
            INIT_RAM_1B => X"003C6666663C000000666666663E000000C6D6FEFE660000003C18181818181C",
            INIT_RAM_1C => X"003E603C067C0000001E0CCCDC760000F0607C6666DC00001E0C7CCCCC760000",
            INIT_RAM_1D => X"006CFEFED6C6000000183C666666000000DC66666666000000305818187C1810",
            INIT_RAM_1E => X"007018180E181870007E4C18327E00003E607C666666000000C66C386CC60000",
            INIT_RAM_1F => X"000000000000000000000000000076DC000E18187018180E0030303000303030"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

end Behavioral; --Gowin_pROM
