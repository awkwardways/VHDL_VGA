//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Sat Aug 23 21:00:56 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [30:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[12:0]})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h60F0F060000000000000A0A00000000040004040000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000402000000000D0E0B0C000000000904020900000000040E0E04000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h40E0400000000000A040E0400000000040202040000000002040402000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h4040202000000000400000000000000000E00000000000002060000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'hE02060E000000000E0C020E000000000E04040C000000000E0A0A0E000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h404020E000000000E0E080C000000000E020C0E00000000020E0A0A000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h206000400000000040004000000000006020E0E000000000E0A0E06000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h400060E0000000004020400000000000E000E000000000002040200000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'hE080806000000000E0A0E0C000000000A0E0A06000000000F05090F000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'hE0A08060000000008080C0E000000000E080C0E000000000C0A0A0C000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'hA0C0C0A000000000E0A0206000000000E04040E000000000A0E0A0A000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'hE0A0A0E000000000A0A0A0E000000000A0E0E0E000000000E080808000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'hE06080E000000000A0C0A0E000000000F0E0A0E00000000080E0A0E000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'hE0E0E0A00000000080C0A0A000000000E0A0A0A000000000404040E000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h6040406000000000E04020E0000000004040E0A000000000A0A040A000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'hF0000000000000000000A0400000000060202060000000002020404000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'hE080600000000000E0A0E08000000000E0E06000000000000000408000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'hC020E0600000000040E0406000000000C0E0E00000000000E0A0E02000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'hA0C0A08000000000C0400040000000004040004000000000A0A0E08000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'hE0A0E00000000000A0A0E00000000000A0E0E00000000000604040C000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'hC0406000000000008080E000000000002060A0400000000080C0A04000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'hE0E0A0000000000040E0A00000000000E0A0A000000000006040604000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h6040C060000000006040C00000000000C060A00000000000A040A00000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h00000000000000000080E02000000000C04060C0000000004040404000000000;

endmodule //Gowin_pROM
