library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity vga_tb is
end entity vga_tb;

architecture sim of vga_tb is 

  constant DATA_BUS_WIDTH    : integer := 16;
  constant SCREEN_WIDTH      : integer := 640;
  constant SCREEN_HEIGHT     : integer := 480;
  constant PX_RESTART_COUNT  : integer := 800;
  constant LN_RESTART_COUNT  : integer := 525;
  constant PX_COUNT_LENGTH   : integer := integer(ceil(log2(real(PX_RESTART_COUNT))));
  constant LN_COUNT_LENGTH   : integer := integer(ceil(log2(real(LN_RESTART_COUNT))));
  constant HS_VISIBLE_AREA   : integer := SCREEN_WIDTH;
  constant HS_FRONT_PORCH    : integer := 16;
  constant HS_SYNC_PULSE     : integer := 96;
  constant HS_BACK_PORCH     : integer := 48;
  constant VS_VISIBLE_AREA   : integer := SCREEN_HEIGHT;
  constant VS_FRONT_PORCH    : integer := 10;
  constant VS_SYNC_PULSE     : integer := 2;
  constant VS_BACK_PORCH     : integer := 33;
  constant ADDRESS_BUS_WIDTH : integer := 15;
  constant VGA_CLK_FREQUENCY : integer := 25e6;
  constant VGA_CLK_PERIOD    : time := 1000 ms / VGA_CLK_FREQUENCY;
  
  signal vga_clk   : std_logic := '1';
  signal ln_enable : std_logic;  
  signal px_count  : std_logic_vector(PX_COUNT_LENGTH - 1 downto 0);
  signal ln_count  : std_logic_vector(LN_COUNT_LENGTH - 1 downto 0);
  signal data_bus  : std_logic_vector(DATA_BUS_WIDTH - 1 downto 0);
  signal hsync     : std_logic;
  signal vsync     : std_logic;
  signal r         : std_logic_vector(4 downto 0);
  signal g         : std_logic_vector(5 downto 0);
  signal b         : std_logic_vector(4 downto 0);
  signal h_visible : std_logic;
  signal v_visible : std_logic;

begin

  
  r <= data_bus(DATA_BUS_WIDTH - 1 downto 11) and (h_visible and v_visible);
  g <= data_bus(10 downto 5) and (h_visible and v_visible);
  b <= data_bus(4 downto 0) and (h_visible and v_visible);
  
  vga_clk <= not vga_clk after VGA_CLK_PERIOD / 2;

  pixelcounter: entity work.px_counter(behavioural)
  generic map (
    RESTART_COUNT => PX_RESTART_COUNT,
    PX_COUNT_LENGTH => PX_COUNT_LENGTH
  )
  port map (
    clk_in => vga_clk,
    px_count => px_count
  );

  linecounter: entity work.ln_counter(behavioural)
  generic map (
    LN_RESTART_COUNT => LN_RESTART_COUNT,
    PX_RESTART_COUNT => PX_RESTART_COUNT,
    PX_COUNT_LENGTH => PX_COUNT_LENGTH,
    LN_COUNT_LENGTH => LN_COUNT_LENGTH
  )
  port map (
    clk_in => vga_clk,
    ln_count => ln_count,
    px_count => px_count
  );

  hsyncgenerator: entity work.hsync_generator(behavioural)
  generic map (
    PX_COUNT_LENGTH => PX_COUNT_LENGTH,
    VISIBLE_AREA => HS_VISIBLE_AREA,
    FRONT_PORCH => HS_FRONT_PORCH,
    SYNC_PULSE => HS_SYNC_PULSE,
    BACK_PORCH => HS_BACK_PORCH 
  )
  port map (
    px_count => px_count, 
    hsync => hsync,
    h_visible => h_visible
  );

  vsyncgenerator: entity work.vsync_generator(behavioural)
  generic map (
    LN_COUNT_LENGTH => LN_COUNT_LENGTH,
    VISIBLE_AREA => VS_VISIBLE_AREA,
    FRONT_PORCH => VS_FRONT_PORCH,
    SYNC_PULSE => VS_SYNC_PULSE,
    BACK_PORCH => VS_BACK_PORCH
  )
  port map (
    vsync => vsync,
    ln_count => ln_count,
    v_visible => v_visible
  );

  rom: entity work.rom(rtl)
  generic map (
    ADDRESS_BUS_WIDTH => ADDRESS_BUS_WIDTH,
    DATA_BUS_WIDTH => DATA_BUS_WIDTH,
    ROM_IMAGE => "scripts\\rom.img"
  )
  port map (
    address_bus => ln_count(6 downto 0) & px_count(7 downto 0),
    data_bus => data_bus,
    chip_select => (h_visible and v_visible),
    clock_in => vga_clk
  ); 
end architecture;